//--------------------------------------------------------------------------//
// Title:        de0_nano_soc_baseline.v                                       //
// Rev:          Rev 0.1                                                    //
// Last Revised: 09/14/2015                                                 //
//--------------------------------------------------------------------------//
// Description: Baseline design file contains DE0 Nano SoC    				 //
//              Board pins and I/O Standards.                               //
//--------------------------------------------------------------------------//
//Copyright 2015 Altera Corporation. All rights reserved.  Altera products
//are protected under numerous U.S. and foreign patents, maskwork rights,
//copyrights and other intellectual property laws.
//                 
//This reference design file, and your use thereof, is subject to and
//governed by the terms and conditions of the applicable Altera Reference
//Design License Agreement.  By using this reference design file, you
//indicate your acceptance of such terms and conditions between you and
//Altera Corporation.  In the event that you do not agree with such terms and
//conditions, you may not use the reference design file. Please promptly                         
//destroy any copies you have made.
//
//This reference design file being provided on an "as-is" basis and as an
//accommodation and therefore all warranties, representations or guarantees
//of any kind (whether express, implied or statutory) including, without
//limitation, warranties of merchantability, non-infringement, or fitness for
//a particular purpose, are specifically disclaimed.  By making this
//reference design file available, Altera expressly does not recommend,
//suggest or require that this reference design file be used in combination 
//with any other product not provided by Altera
//----------------------------------------------------------------------------

//Group Enable Definitions
//This lists every pinout group
//Users can enable any group by uncommenting the corresponding line below:
//`define enable_ADC
//`define enable_ARDUINO
//`define enable_GPIO0
//`define enable_GPIO1
//`define enable_HPS

module proj_agh(


	//////////// CLOCK //////////
	input 		          		FPGA_CLK_50,
	input 		          		FPGA_CLK2_50,
	input 		          		FPGA_CLK3_50,

`ifdef enable_ADC
	//////////// ADC //////////
	/* 3.3-V LVTTL */
	output		          		ADC_CONVST,
	output		          		ADC_SCLK,
	output		          		ADC_SDI,
	input 		          		ADC_SDO,
`endif
	
`ifdef enable_ARDUINO
	//////////// ARDUINO ////////////
	/* 3.3-V LVTTL */
	inout					[15:0]	ARDUINO_IO,
	inout								ARDUINO_RESET_N,
`endif
	
`ifdef enable_GPIO0
	//////////// GPIO 0 ////////////
	/* 3.3-V LVTTL */
	inout				[35:0]		GPIO_0,
`endif

`ifdef enable_GPIO1	
	//////////// GPIO 1 ////////////
	/* 3.3-V LVTTL */
	inout				[35:0]		GPIO_1,
`endif

`ifdef enable_HPS
	//////////// HPS //////////
	/* 3.3-V LVTTL */
	inout 		          		HPS_CONV_USB_N,
	
	/* SSTL-15 Class I */
	output		    [14:0]		HPS_DDR3_ADDR,
	output		     [2:0]		HPS_DDR3_BA,
	output		          		HPS_DDR3_CAS_N,
	output		          		HPS_DDR3_CKE,
	output		          		HPS_DDR3_CS_N,
	output		     [3:0]		HPS_DDR3_DM,
	inout 		    [31:0]		HPS_DDR3_DQ,
	output		          		HPS_DDR3_ODT,
	output		          		HPS_DDR3_RAS_N,
	output		          		HPS_DDR3_RESET_N,
	input 		          		HPS_DDR3_RZQ,
	output		          		HPS_DDR3_WE_N,
	/* DIFFERENTIAL 1.5-V SSTL CLASS I */
	output		          		HPS_DDR3_CK_N,
	output		          		HPS_DDR3_CK_P,
	inout 		     [3:0]		HPS_DDR3_DQS_N,
	inout 		     [3:0]		HPS_DDR3_DQS_P,
	
	/* 3.3-V LVTTL */
	output		          		HPS_ENET_GTX_CLK,
	inout 		          		HPS_ENET_INT_N,
	output		          		HPS_ENET_MDC,
	inout 		          		HPS_ENET_MDIO,
	input 		          		HPS_ENET_RX_CLK,
	input 		     [3:0]		HPS_ENET_RX_DATA,
	input 		          		HPS_ENET_RX_DV,
	output		     [3:0]		HPS_ENET_TX_DATA,
	output		          		HPS_ENET_TX_EN,
	inout 		          		HPS_GSENSOR_INT,
	inout 		          		HPS_I2C0_SCLK,
	inout 		          		HPS_I2C0_SDAT,
	inout 		          		HPS_I2C1_SCLK,
	inout 		          		HPS_I2C1_SDAT,
	inout 		          		HPS_KEY,
	inout 		          		HPS_LED,
	inout 		          		HPS_LTC_GPIO,
	output		          		HPS_SD_CLK,
	inout 		          		HPS_SD_CMD,
	inout 		     [3:0]		HPS_SD_DATA,
	output		          		HPS_SPIM_CLK,
	input 		          		HPS_SPIM_MISO,
	output		          		HPS_SPIM_MOSI,
	inout 		          		HPS_SPIM_SS,
	input 		          		HPS_UART_RX,
	output		          		HPS_UART_TX,
	input 		          		HPS_USB_CLKOUT,
	inout 		     [7:0]		HPS_USB_DATA,
	input 		          		HPS_USB_DIR,
	input 		          		HPS_USB_NXT,
	output		          		HPS_USB_STP,
`endif
	
	//////////// KEY ////////////
	/* 3.3-V LVTTL */
	input				[1:0]			KEY,
	
	//////////// LED ////////////
	/* 3.3-V LVTTL */
	//output			[7:0]			LED,
	
	//////////// SW ////////////
	/* 3.3-V LVTTL */
	input				[3:0]			SW

);


localparam WIDTH = 32;

wire rst;
wire pll_rst;
wire pll_clk;
wire pll_lock;

wire [WIDTH-1:0]		alu_data_a;
wire [WIDTH-1:0]		alu_data_b;
wire [(WIDTH*2)-1:0]	alu_out;
wire [7:0] 				alu_ops;

wire [4:0]	rom_addr;
wire 		rom_clk;
wire 		rom_rd;
wire [31:0] rom_data;

wire [4:0]	mem_a_addr;
wire 		mem_a_clk;
wire [31:0]	mem_a_wrdata;
wire 		mem_a_rd;
wire 		mem_a_wr;
wire [31:0]	mem_a_data;

wire [4:0]	mem_b_addr;
wire 		mem_b_clk;
wire [31:0]	mem_b_wrdata;
wire 		mem_b_rd;
wire 		mem_b_wr;
wire [31:0]	mem_b_data;

wire [4:0]	mem_c_addr;
wire 		mem_c_clk;
wire [63:0]	mem_c_wrdata;
wire 		mem_c_rd;
wire 		mem_c_wr;
wire [63:0]	mem_c_data;


//--- RTL ---


power_ctrl INST_POWER_CTRL(

    .ref_clk	(FPGA_CLK_50)
    ,.ref_rst	(KEY)

    ,.rom_clk	(rom_clk)
    ,.mem_a_clk	(mem_a_clk)
    ,.mem_b_clk	(mem_b_clk)
    ,.mem_c_clk	(mem_c_clk)
    ,.ctrl_clk	(ctrl_clk)
    ,.rst		(rst)
);


//assign rom_clk = pll_clk;

gen_rom	INST_ROM (
	.address	( rom_addr )
	,.clock 	( rom_clk )
	,.rden		( rom_rd )
	,.q			( rom_data )
	);



//assign mem_a_clk = pll_clk;

gen_ram	INST_RAM_DATA_A (
	 .address ( mem_a_addr )
	,.clock   ( mem_a_clk )
	,.data    ( mem_a_wrdata )
	,.rden    ( mem_a_rd )
	,.wren    ( )
	,.q       ( mem_a_data )
	);



//assign mem_b_clk = pll_clk;

gen_ram	INST_RAM_DATA_B (
	 .address ( mem_b_addr )
	,.clock   ( mem_b_clk )
	,.data    ( mem_b_wrdata )
	,.rden    ( mem_b_rd )
	,.wren    ( )
	,.q       ( mem_b_data )
	);



//assign mem_c_clk = pll_clk;

assign mem_c_wrdata = alu_out;

gen_ram_C	INST_RAM_DATA_C (
	 .address ( mem_c_addr )
	,.clock   ( mem_c_clk )
	,.data    ( mem_c_wrdata )
//	,.rden    ( mem_c_rd )
	,.wren    ( mem_c_wr)
	,.q       ( mem_c_data )
	);




assign GPIO_0		= {4'h0, alu_out[31:0]};
assign alu_data_a	= mem_a_data;
assign alu_data_b	= mem_b_data;


alu 
	#(
		.WIDTH (WIDTH) 
	)
	INST_ALU
	(
	 .inputA	(alu_data_a)
	,.inputB	(alu_data_b)
	,.operation	(alu_ops)
	
	,.outputC	(alu_out)

	);



ctrl INST_CTRL(
    .clk			(ctrl_clk)
    ,.rst			(rst)

    ,.rom_addr		(rom_addr)
    ,.rom_rd		(rom_rd)
    ,.rom_data		(rom_data)

    ,.mem_a_rd		(mem_a_rd)
    ,.mem_a_addr	(mem_a_addr)
    ,.mem_b_rd		(mem_b_rd)
    ,.mem_b_addr	(mem_b_addr)
    ,.mem_c_wr		(mem_c_wr)
    ,.mem_c_addr	(mem_c_addr)

    ,.ops			(alu_ops)

);



endmodule
